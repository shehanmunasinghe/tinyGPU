module control_unit (
    ports //TODO
);
    
endmodule