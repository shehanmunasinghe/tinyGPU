/*************************************************
        Make a copy of this file and name it as 'constants_local.v', edit the filepaths accodingly
*************************************************/

//To know whether constants has been included. If not will use local definitions inside modules.
`define INC_CONSTANTS_LOCAL 1

/*************************************************
    Local Constants - eg: memory file paths, etc
    This will not be tracked by git
*************************************************/

// Instruction memory
`define INSTMEM_FILEPATH "PleaseSpecifyAFilePath"

//Data memory
`define DATAMEM_FILEPATH "PleaseSpecifyAFilePath"