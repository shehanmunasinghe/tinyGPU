module scheduler (
    ports //TODO
);
    
endmodule